netcdf std14profile {
dimensions:
	time = 1, depth = 31, lat = 30, lon = 30;
variables:
	float time(time), depth(depth), lat(lat), lon(lon), speed(time,depth,lat,lon);
	depth:units = "meters";
	lat:units = "degrees_north";
	lon:units = "degrees_east";
	speed:units = "meters/sec";
data:
	time = 0 ;
	depth = -0.000,-10.000,-20.000,-30.000,-50.000,-75.000,-100.000,-125.000,-150.000,-200.000,-250.000,-300.000,-400.000,-500.000,-600.000,-700.000,-800.000,-900.000,-1000.000,-1100.000,-1200.000,-1300.000,-1400.000,-1500.000,-1750.000,-2000.000,-2500.000,-3000.000,-4000.000,-5000.000,-5530;
	lat = 16.123,16.418,16.714,17.010,17.305,17.601,17.897,18.193,18.488,18.784,19.080,19.375,19.671,19.967,20.262,20.558,20.854,21.150,21.445,21.741,22.037,22.332,22.628,22.924,23.220,23.515,23.811,24.107,24.402,2.469805e+001;
	lon = -164.654,-164.341,-164.027,-163.713,-163.400,-163.086,-162.772,-162.459,-162.145,-161.831,-161.518,-161.204,-160.890,-160.577,-160.263,-159.949,-159.636,-159.322,-159.008,-158.695,-158.381,-158.067,-157.754,-157.440,-157.126,-156.813,-156.499,-156.185,-155.872,-1.555578e+002;
	speed = 
		1534.64,1534.64,1534.41,1534.21,1534.21,1534.13,1534.13,1534.04,1533.99,1533.99,1533.93,1533.85,1533.85,1533.78,1533.78,1533.73,1533.67,1533.67,1533.51,1533.29,1533.29,1533.29,1533.29,1533.29,1533.29,1533.29,1533.29,1533.29,1533.29,1533.29,
		1534.63,1534.63,1534.38,1534.23,1534.23,1534.06,1534.06,1533.96,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,
		1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,
		1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,
		1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,
		1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,
		1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,
		1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,
		1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,
		1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,
		1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,
		1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,
		1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,
		1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,
		1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,
		1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,
		1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,
		1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,
		1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,
		1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,
		1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,
		1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,
		1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,
		1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,
		1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,
		1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,
		1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,
		1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,
		1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,
		1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,1533.89,
		
		1534.79,1534.79,1534.58,1534.38,1534.38,1534.29,1534.29,1534.21,1534.16,1534.16,1534.10,1534.02,1534.02,1533.95,1533.95,1533.90,1533.84,1533.84,1533.68,1533.46,1533.46,1533.46,1533.46,1533.46,1533.46,1533.46,1533.46,1533.46,1533.46,1533.46,
		1534.79,1534.79,1534.55,1534.39,1534.39,1534.23,1534.23,1534.12,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,
		1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,
		1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,
		1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,
		1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,
		1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,
		1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,
		1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,
		1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,
		1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,
		1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,
		1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,
		1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,
		1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,
		1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,
		1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,
		1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,
		1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,
		1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,
		1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,
		1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,
		1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,
		1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,
		1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,
		1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,
		1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,
		1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,
		1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,
		1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,1534.06,
		
		1534.96,1534.96,1534.74,1534.55,1534.55,1534.45,1534.45,1534.37,1534.32,1534.32,1534.26,1534.18,1534.18,1534.11,1534.11,1534.07,1533.99,1533.99,1533.84,1533.62,1533.62,1533.62,1533.62,1533.62,1533.62,1533.62,1533.62,1533.62,1533.62,1533.62,
		1534.96,1534.96,1534.71,1534.54,1534.54,1534.40,1534.40,1534.29,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,
		1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,
		1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,
		1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,
		1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,
		1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,
		1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,
		1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,
		1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,
		1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,
		1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,
		1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,
		1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,
		1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,
		1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,
		1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,
		1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,
		1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,
		1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,
		1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,
		1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,
		1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,
		1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,
		1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,
		1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,
		1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,
		1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,
		1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,
		1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,1534.22,
		
		1535.15,1535.15,1534.93,1534.73,1534.73,1534.59,1534.59,1534.55,1534.49,1534.49,1534.43,1534.35,1534.35,1534.28,1534.28,1534.23,1534.17,1534.17,1534.01,1533.79,1533.79,1533.79,1533.79,1533.79,1533.79,1533.79,1533.79,1533.79,1533.79,1533.79,
		1535.14,1535.14,1534.90,1534.73,1534.73,1534.57,1534.57,1534.46,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,
		1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,
		1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,
		1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,
		1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,
		1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,
		1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,
		1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,
		1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,
		1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,
		1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,
		1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,
		1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,
		1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,
		1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,
		1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,
		1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,
		1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,
		1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,
		1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,
		1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,
		1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,
		1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,
		1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,
		1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,
		1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,
		1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,
		1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,
		1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,1534.39,
		
		1535.50,1535.50,1535.26,1535.10,1535.10,1534.92,1534.92,1534.82,1534.81,1534.81,1534.73,1534.65,1534.65,1534.56,1534.56,1534.51,1534.41,1534.41,1534.28,1534.03,1534.03,1534.03,1534.03,1534.03,1534.03,1534.03,1534.03,1534.03,1534.03,1534.03,
		1535.53,1535.53,1535.30,1535.07,1535.07,1534.91,1534.91,1534.79,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		
		1535.65,1535.65,1535.38,1535.27,1535.27,1534.90,1534.90,1534.78,1534.95,1534.95,1534.85,1534.73,1534.73,1534.56,1534.56,1534.58,1534.32,1534.32,1534.20,1533.92,1533.92,1533.92,1533.92,1533.92,1533.92,1533.92,1533.92,1533.92,1533.92,1533.92,
		1535.89,1535.89,1535.52,1535.21,1535.21,1535.00,1535.00,1534.88,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,1534.69,
		
		1534.88,1534.88,1534.51,1534.46,1534.46,1533.76,1533.76,1533.62,1534.04,1534.04,1533.92,1533.78,1533.78,1533.55,1533.55,1533.65,1533.18,1533.18,1532.93,1532.52,1532.52,1532.52,1532.52,1532.52,1532.52,1532.52,1532.52,1532.52,1532.52,1532.52,
		1535.63,1535.63,1535.02,1534.51,1534.51,1534.16,1534.16,1533.99,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,
		1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,
		1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,
		1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,
		1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,
		1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,
		1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,
		1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,
		1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,
		1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,
		1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,
		1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,
		1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,
		1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,
		1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,
		1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,
		1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,
		1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,
		1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,
		1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,
		1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,
		1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,
		1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,
		1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,
		1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,
		1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,
		1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,
		1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,
		1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,1533.69,
		
		1532.52,1532.52,1531.94,1531.74,1531.74,1530.75,1530.75,1530.49,1531.16,1531.16,1530.94,1530.96,1530.96,1530.64,1530.64,1530.90,1530.19,1530.19,1529.76,1529.11,1529.11,1529.11,1529.11,1529.11,1529.11,1529.11,1529.11,1529.11,1529.11,1529.11,
		1534.16,1534.16,1533.04,1532.14,1532.14,1531.65,1531.65,1531.35,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,
		1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,
		1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,
		1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,
		1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,
		1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,
		1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,
		1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,
		1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,
		1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,
		1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,
		1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,
		1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,
		1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,
		1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,
		1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,
		1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,
		1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,
		1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,
		1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,
		1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,
		1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,
		1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,
		1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,
		1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,
		1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,
		1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,
		1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,
		1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,1531.01,
		
		1527.94,1527.94,1527.16,1526.57,1526.57,1525.65,1525.65,1525.13,1525.75,1525.75,1525.39,1525.73,1525.73,1525.45,1525.45,1525.81,1525.13,1525.13,1524.46,1523.55,1523.55,1523.55,1523.55,1523.55,1523.55,1523.55,1523.55,1523.55,1523.55,1523.55,
		1530.71,1530.71,1528.99,1527.67,1527.67,1527.02,1527.02,1526.56,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,
		1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,
		1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,
		1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,
		1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,
		1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,
		1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,
		1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,
		1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,
		1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,
		1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,
		1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,
		1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,
		1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,
		1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,
		1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,
		1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,
		1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,
		1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,
		1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,
		1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,
		1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,
		1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,
		1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,
		1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,
		1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,
		1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,
		1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,
		1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,1526.28,
		
		1514.21,1514.21,1513.39,1512.15,1512.15,1512.05,1512.05,1511.33,1511.28,1511.28,1510.96,1511.74,1511.74,1511.77,1511.77,1512.15,1511.96,1511.96,1511.13,1510.24,1510.24,1510.24,1510.24,1510.24,1510.24,1510.24,1510.24,1510.24,1510.24,1510.24,
		1518.06,1518.06,1515.77,1514.45,1514.45,1513.76,1513.76,1513.27,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,
		1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,
		1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,
		1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,
		1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,
		1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,
		1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,
		1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,
		1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,
		1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,
		1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,
		1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,
		1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,
		1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,
		1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,
		1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,
		1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,
		1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,
		1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,
		1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,
		1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,
		1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,
		1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,
		1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,
		1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,
		1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,
		1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,
		1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,
		1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,1513.42,
		
		1502.30,1502.30,1501.77,1501.64,1501.64,1501.13,1501.13,1501.03,1501.16,1501.16,1501.43,1501.74,1501.74,1501.75,1501.75,1502.24,1501.80,1501.80,1501.31,1500.72,1500.72,1500.72,1500.72,1500.72,1500.72,1500.72,1500.72,1500.72,1500.72,1500.72,
		1505.52,1505.52,1503.65,1502.98,1502.98,1502.74,1502.74,1502.81,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,
		1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,
		1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,
		1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,
		1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,
		1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,
		1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,
		1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,
		1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,
		1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,
		1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,
		1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,
		1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,
		1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,
		1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,
		1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,
		1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,
		1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,
		1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,
		1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,
		1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,
		1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,
		1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,
		1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,
		1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,
		1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,
		1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,
		1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,
		1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,1502.84,
		
		1496.23,1496.23,1495.84,1496.52,1496.52,1496.10,1496.10,1496.02,1496.75,1496.75,1496.63,1497.05,1497.05,1497.06,1497.06,1497.50,1497.14,1497.14,1497.01,1496.78,1496.78,1496.78,1496.78,1496.78,1496.78,1496.78,1496.78,1496.78,1496.78,1496.78,
		1498.53,1498.53,1497.37,1496.94,1496.94,1497.03,1497.03,1497.36,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,
		1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,
		1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,
		1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,
		1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,
		1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,
		1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,
		1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,
		1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,
		1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,
		1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,
		1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,
		1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,
		1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,
		1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,
		1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,
		1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,
		1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,
		1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,
		1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,
		1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,
		1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,
		1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,
		1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,
		1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,
		1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,
		1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,
		1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,
		1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,1497.15,
		
		1488.02,1488.02,1488.49,1488.80,1488.80,1488.75,1488.75,1488.59,1488.60,1488.60,1488.82,1489.58,1489.58,1490.11,1490.11,1490.59,1490.93,1490.93,1491.13,1491.52,1491.52,1491.52,1491.52,1491.52,1491.52,1491.52,1491.52,1491.52,1491.52,1491.52,
		1488.44,1488.44,1488.60,1488.94,1488.94,1488.93,1488.93,1488.74,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,
		1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,
		1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,
		1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,
		1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,
		1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,
		1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,
		1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,
		1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,
		1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,
		1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,
		1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,
		1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,
		1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,
		1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,
		1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,
		1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,
		1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,
		1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,
		1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,
		1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,
		1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,
		1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,
		1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,
		1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,
		1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,
		1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,
		1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,
		1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,1488.72,
		
		1484.97,1484.97,1485.20,1485.24,1485.24,1485.18,1485.18,1485.11,1485.17,1485.17,1485.50,1486.28,1486.28,1486.68,1486.68,1487.06,1487.52,1487.52,1487.80,1488.49,1488.49,1488.49,1488.49,1488.49,1488.49,1488.49,1488.49,1488.49,1488.49,1488.49,
		1484.93,1484.93,1484.92,1485.01,1485.01,1484.94,1484.94,1484.84,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,
		1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,
		1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,
		1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,
		1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,
		1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,
		1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,
		1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,
		1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,
		1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,
		1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,
		1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,
		1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,
		1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,
		1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,
		1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,
		1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,
		1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,
		1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,
		1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,
		1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,
		1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,
		1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,
		1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,
		1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,
		1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,
		1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,
		1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,
		1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,
		
		1484.77,1484.77,1484.65,1484.55,1484.55,1484.59,1484.59,1484.63,1484.83,1484.83,1485.12,1485.53,1485.53,1485.49,1485.49,1485.50,1485.87,1485.87,1486.22,1486.85,1486.85,1486.85,1486.85,1486.85,1486.85,1486.85,1486.85,1486.85,1486.85,1486.85,
		1484.52,1484.52,1484.36,1484.28,1484.28,1484.20,1484.20,1484.28,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,
		1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,
		1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,
		1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,
		1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,
		1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,
		1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,
		1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,
		1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,
		1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,
		1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,
		1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,
		1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,
		1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,
		1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,
		1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,
		1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,
		1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,
		1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,
		1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,
		1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,
		1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,
		1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,
		1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,
		1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,
		1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,
		1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,
		1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,
		1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,1484.46,
		
		1484.37,1484.37,1484.33,1484.37,1484.37,1484.53,1484.53,1484.85,1485.05,1485.05,1485.17,1485.39,1485.39,1485.24,1485.24,1485.08,1485.35,1485.35,1485.59,1486.15,1486.15,1486.15,1486.15,1486.15,1486.15,1486.15,1486.15,1486.15,1486.15,1486.15,
		1484.14,1484.14,1484.06,1484.11,1484.11,1484.19,1484.19,1484.40,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		
		1484.34,1484.34,1484.32,1484.41,1484.41,1484.61,1484.61,1484.93,1485.14,1485.14,1485.23,1485.28,1485.28,1485.08,1485.08,1484.92,1485.03,1485.03,1485.23,1485.63,1485.63,1485.63,1485.63,1485.63,1485.63,1485.63,1485.63,1485.63,1485.63,1485.63,
		1484.12,1484.12,1484.05,1484.10,1484.10,1484.22,1484.22,1484.50,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,
		1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,
		1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,
		1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,
		1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,
		1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,
		1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,
		1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,
		1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,
		1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,
		1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,
		1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,
		1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,
		1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,
		1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,
		1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,
		1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,
		1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,
		1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,
		1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,
		1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,
		1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,
		1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,
		1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,
		1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,
		1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,
		1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,
		1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,
		1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,1484.69,
		
		1484.35,1484.35,1484.31,1484.35,1484.35,1484.55,1484.55,1484.76,1484.92,1484.92,1484.97,1484.97,1484.97,1484.77,1484.77,1484.59,1484.66,1484.66,1484.81,1485.11,1485.11,1485.11,1485.11,1485.11,1485.11,1485.11,1485.11,1485.11,1485.11,1485.11,
		1484.18,1484.18,1484.10,1484.10,1484.10,1484.18,1484.18,1484.39,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,1484.52,
		
		1484.34,1484.34,1484.30,1484.30,1484.30,1484.27,1484.27,1484.42,1484.51,1484.51,1484.51,1484.55,1484.55,1484.38,1484.38,1484.27,1484.40,1484.40,1484.52,1484.68,1484.68,1484.68,1484.68,1484.68,1484.68,1484.68,1484.68,1484.68,1484.68,1484.68,
		1484.26,1484.26,1484.18,1484.09,1484.09,1484.09,1484.09,1484.13,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,
		1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,
		1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,
		1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,
		1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,
		1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,
		1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,
		1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,
		1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,
		1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,
		1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,
		1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,
		1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,
		1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,
		1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,
		1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,
		1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,
		1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,
		1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,
		1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,
		1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,
		1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,
		1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,
		1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,
		1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,
		1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,
		1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,
		1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,
		1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,1484.18,
		
		1484.49,1484.49,1484.39,1484.27,1484.27,1484.22,1484.22,1484.20,1484.20,1484.20,1484.18,1484.21,1484.21,1484.17,1484.17,1484.13,1484.28,1484.28,1484.42,1484.68,1484.68,1484.68,1484.68,1484.68,1484.68,1484.68,1484.68,1484.68,1484.68,1484.68,
		1484.41,1484.41,1484.28,1484.15,1484.15,1483.99,1483.99,1483.99,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,
		1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,
		1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,
		1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,
		1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,
		1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,
		1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,
		1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,
		1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,
		1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,
		1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,
		1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,
		1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,
		1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,
		1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,
		1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,
		1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,
		1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,
		1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,
		1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,
		1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,
		1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,
		1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,
		1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,
		1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,
		1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,
		1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,
		1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,
		1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,1483.94,
		
		1484.81,1484.81,1484.68,1484.47,1484.47,1484.39,1484.39,1484.26,1484.22,1484.22,1484.18,1484.29,1484.29,1484.25,1484.25,1484.28,1484.48,1484.48,1484.69,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,1484.93,
		1484.74,1484.74,1484.56,1484.39,1484.39,1484.23,1484.23,1484.09,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,
		1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,
		1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,
		1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,
		1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,
		1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,
		1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,
		1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,
		1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,
		1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,
		1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,
		1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,
		1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,
		1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,
		1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,
		1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,
		1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,
		1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,
		1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,
		1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,
		1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,
		1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,
		1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,
		1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,
		1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,
		1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,
		1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,
		1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,
		1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,1484.01,
		
		1485.34,1485.34,1485.21,1485.04,1485.04,1484.87,1484.87,1484.74,1484.61,1484.61,1484.61,1484.77,1484.77,1484.77,1484.77,1484.84,1485.00,1485.00,1485.26,1485.54,1485.54,1485.54,1485.54,1485.54,1485.54,1485.54,1485.54,1485.54,1485.54,1485.54,
		1485.31,1485.31,1485.04,1484.95,1484.95,1484.74,1484.74,1484.57,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,
		1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,
		1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,
		1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,
		1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,
		1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,
		1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,
		1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,
		1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,
		1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,
		1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,
		1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,
		1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,
		1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,
		1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,
		1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,
		1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,
		1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,
		1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,
		1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,
		1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,
		1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,
		1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,
		1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,
		1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,
		1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,
		1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,
		1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,
		1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,1484.48,
		
		1486.12,1486.12,1485.99,1485.76,1485.76,1485.72,1485.72,1485.63,1485.55,1485.55,1485.55,1485.58,1485.58,1485.62,1485.62,1485.70,1485.88,1485.88,1486.08,1486.38,1486.38,1486.38,1486.38,1486.38,1486.38,1486.38,1486.38,1486.38,1486.38,1486.38,
		1486.07,1486.07,1485.90,1485.73,1485.73,1485.59,1485.59,1485.46,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,
		1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,
		1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,
		1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,
		1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,
		1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,
		1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,
		1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,
		1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,
		1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,
		1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,
		1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,
		1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,
		1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,
		1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,
		1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,
		1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,
		1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,
		1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,
		1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,
		1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,
		1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,
		1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,
		1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,
		1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,
		1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,
		1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,
		1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,
		1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,1485.33,
		
		1487.01,1487.01,1486.92,1486.84,1486.84,1486.74,1486.74,1486.70,1486.70,1486.70,1486.65,1486.74,1486.74,1486.70,1486.70,1486.73,1486.90,1486.90,1487.03,1487.38,1487.38,1487.38,1487.38,1487.38,1487.38,1487.38,1487.38,1487.38,1487.38,1487.38,
		1487.01,1487.01,1486.84,1486.75,1486.75,1486.65,1486.65,1486.57,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,
		1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,
		1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,
		1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,
		1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,
		1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,
		1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,
		1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,
		1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,
		1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,
		1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,
		1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,
		1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,
		1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,
		1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,
		1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,
		1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,
		1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,
		1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,
		1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,
		1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,
		1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,
		1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,
		1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,
		1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,
		1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,
		1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,
		1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,
		1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,1486.48,
		
		1489.50,1489.50,1489.45,1489.45,1489.45,1489.50,1489.50,1489.54,1489.57,1489.57,1489.53,1489.53,1489.53,1489.44,1489.44,1489.35,1489.50,1489.50,1489.54,1489.71,1489.71,1489.71,1489.71,1489.71,1489.71,1489.71,1489.71,1489.71,1489.71,1489.71,
		1489.50,1489.50,1489.45,1489.37,1489.37,1489.37,1489.37,1489.44,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,
		1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,
		1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,
		1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,
		1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,
		1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,
		1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,
		1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,
		1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,
		1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,
		1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,
		1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,
		1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,
		1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,
		1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,
		1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,
		1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,
		1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,
		1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,
		1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,
		1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,
		1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,
		1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,
		1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,
		1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,
		1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,
		1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,
		1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,
		1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,1489.48,
		
		1492.40,1492.40,1492.44,1492.46,1492.46,1492.53,1492.53,1492.62,1492.68,1492.68,1492.64,1492.59,1492.59,1492.46,1492.46,1492.44,1492.40,1492.40,1492.40,1492.50,1492.50,1492.50,1492.50,1492.50,1492.50,1492.50,1492.50,1492.50,1492.50,1492.50,
		1492.37,1492.37,1492.37,1492.42,1492.42,1492.51,1492.51,1492.55,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,
		1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,
		1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,
		1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,
		1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,
		1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,
		1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,
		1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,
		1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,
		1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,
		1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,
		1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,
		1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,
		1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,
		1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,
		1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,
		1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,
		1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,
		1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,
		1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,
		1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,
		1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,
		1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,
		1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,
		1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,
		1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,
		1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,
		1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,
		1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,1492.64,
		
		1499.48,1499.48,1499.52,1499.57,1499.57,1499.61,1499.61,1499.70,1499.70,1499.70,1499.70,1499.70,1499.70,1499.61,1499.61,1499.57,1499.52,1499.52,1499.49,1499.49,1499.49,1499.49,1499.49,1499.49,1499.49,1499.49,1499.49,1499.49,1499.49,1499.49,
		1499.48,1499.48,1499.52,1499.57,1499.57,1499.65,1499.65,1499.70,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,
		1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,
		1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,
		1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,
		1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,
		1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,
		1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,
		1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,
		1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,
		1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,
		1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,
		1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,
		1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,
		1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,
		1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,
		1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,
		1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,
		1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,
		1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,
		1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,
		1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,
		1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,
		1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,
		1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,
		1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,
		1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,
		1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,
		1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,
		1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,1499.68,
		
		1507.51,1507.51,1507.51,1507.51,1507.51,1507.51,1507.51,1507.51,1507.60,1507.60,1507.60,1507.60,1507.60,1507.51,1507.51,1507.51,1507.51,1507.51,1507.51,1507.51,1507.51,1507.51,1507.51,1507.51,1507.51,1507.51,1507.51,1507.51,1507.51,1507.51,
		1507.51,1507.51,1507.51,1507.51,1507.51,1507.51,1507.51,1507.51,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,
		1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,
		1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,
		1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,
		1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,
		1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,
		1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,
		1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,
		1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,
		1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,
		1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,
		1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,
		1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,
		1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,
		1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,
		1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,
		1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,
		1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,
		1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,
		1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,
		1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,
		1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,
		1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,
		1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,
		1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,
		1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,
		1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,
		1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,
		1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,1507.60,
		
		1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,
		1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.50,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,
		1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,
		1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,
		1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,
		1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,
		1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,
		1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,
		1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,
		1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,
		1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,
		1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,
		1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,
		1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,
		1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,
		1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,
		1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,
		1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,
		1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,
		1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,
		1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,
		1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,
		1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,
		1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,
		1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,
		1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,
		1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,
		1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,
		1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,
		1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,1524.41,
		
		1542.39,1542.39,1542.39,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.50,1542.50,1542.50,1542.50,1542.50,1542.50,1542.50,1542.50,1542.50,1542.50,1542.50,1542.50,1542.50,1542.50,
		1542.39,1542.39,1542.48,1542.48,1542.48,1542.48,1542.48,1542.52,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,
		1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,
		1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,
		1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,
		1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,
		1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,
		1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,
		1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,
		1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,
		1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,
		1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,
		1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,
		1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,
		1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,
		1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,
		1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,
		1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,
		1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,
		1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,
		1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,
		1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,
		1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,
		1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,
		1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,
		1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,
		1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,
		1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,
		1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,
		1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,1542.48,
		
		1552.49,1552.49,1552.49,1552.40,1552.40,1554.46,1554.46,1554.46,1553.87,1553.87,1553.91,1554.34,1554.34,1554.17,1554.17,1555.68,1554.58,1554.58,1554.60,1558.19,1558.19,1558.19,1558.19,1558.19,1558.19,1558.19,1558.19,1558.19,1558.19,1558.19,
		1552.04,1552.04,1552.76,1553.24,1553.24,1554.07,1554.07,1553.34,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,
		1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,
		1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,
		1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,
		1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,
		1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,
		1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,
		1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,
		1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,
		1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,
		1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,
		1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,
		1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,
		1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,
		1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,
		1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,
		1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,
		1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,
		1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,
		1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,
		1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,
		1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,
		1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,
		1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,
		1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,
		1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,
		1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,
		1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,
		1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17,1554.17
		
			;
}
