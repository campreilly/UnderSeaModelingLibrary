netcdf std14bathy {
dimensions:
	lat = 60, lon = 59;
variables:
	float lat(lat), lon(lon), depth(lat,lon);
	lat:units = "degrees_north";
	lon:units = "degrees_east";
	depth:units = "meters";
data:
	lat = 16.122,16.270,16.418,16.566,16.713,16.861,17.009,17.157,17.305,17.453,17.601,17.748,17.896,18.044,18.192,18.340,18.488,18.636,18.783,18.931,19.079,19.227,19.375,19.523,19.671,19.818,19.966,20.114,20.262,20.410,20.558,20.706,20.853,21.001,21.149,21.297,21.445,21.593,21.740,21.888,22.036,22.184,22.332,22.480,22.628,22.775,22.923,23.071,23.219,23.367,23.515,23.663,23.810,23.958,24.106,24.254,24.402,24.550,24.698,2.484500e+001;
	lon = -164.497,-164.340,-164.183,-164.027,-163.870,-163.713,-163.556,-163.399,-163.242,-163.086,-162.929,-162.772,-162.615,-162.458,-162.301,-162.145,-161.988,-161.831,-161.674,-161.517,-161.360,-161.204,-161.047,-160.890,-160.733,-160.576,-160.419,-160.262,-160.106,-159.949,-159.792,-159.635,-159.478,-159.321,-159.165,-159.008,-158.851,-158.694,-158.537,-158.380,-158.224,-158.067,-157.910,-157.753,-157.596,-157.439,-157.283,-157.126,-156.969,-156.812,-156.655,-156.498,-156.342,-156.185,-156.028,-155.871,-155.714,-155.557,-1.554010e+002;
	depth = 
		-5502,-5514,-5507,-5499,-5508,-5512,-5511,-5500,-5519,-5550,-5576,-5620,-5447,-5327,-4298,-5236,-4966,-3753,-4522,-5006,-5575,-5585,-5593,-5596,-5587,-5554,-5510,-5465,-5429,-5432,-5253,-5513,-5587,-5572,-5529,-5498,-5552,-5600,-5773,-5526,-5393,-5214,-5393,-5395,-5296,-5195,-5190,-5283,-5282,-5223,-5051,-5132,-5137,-5175,-4689,-4754,-4930,-4999,-5059,
		-5495,-5506,-5500,-5505,-5519,-5523,-5503,-5501,-5514,-5508,-5569,-5554,-5478,-5176,-5472,-5458,-3487,-4996,-5334,-5549,-5591,-5598,-5620,-5621,-5612,-5595,-5575,-5572,-5603,-5689,-5597,-5396,-5440,-5451,-5369,-5307,-5340,-5505,-5588,-5585,-5398,-5399,-5406,-5358,-5226,-5125,-4552,-5184,-5119,-5072,-5105,-5104,-5181,-4982,-4071,-4255,-4477,-4985,-5000,
		-5492,-5489,-5500,-5504,-5512,-5514,-5504,-5522,-5517,-5559,-5541,-5446,-4999,-4400,-5466,-5266,-5471,-5481,-5555,-5564,-5598,-5617,-5621,-5619,-5608,-5596,-5593,-5601,-5631,-5707,-5699,-5599,-5410,-5402,-5355,-5239,-5192,-5418,-5413,-5402,-5387,-5399,-5394,-5375,-5243,-5170,-5192,-5064,-5135,-5074,-5125,-5187,-5184,-4913,-4916,-4985,-4988,-4993,-4993,
		-5439,-5478,-5497,-5501,-5529,-5531,-5506,-5559,-5549,-5589,-5540,-4988,-4566,-4400,-5333,-5540,-5528,-5544,-5559,-5585,-5600,-5602,-5602,-5600,-5599,-5599,-5601,-5611,-5627,-5618,-5603,-5563,-5471,-5406,-5389,-5398,-5399,-5400,-5395,-5379,-5307,-5293,-5282,-5206,-5173,-5191,-5194,-5189,-5155,-5117,-5059,-5096,-5100,-4994,-4988,-4987,-4980,-4973,-4952,
		-5474,-5498,-5500,-5502,-5525,-5518,-5523,-5477,-5551,-5609,-5469,-3414,-5009,-5476,-5567,-5603,-5581,-5592,-5597,-5592,-5580,-5569,-5569,-5572,-5585,-5603,-5605,-5606,-5612,-5635,-5630,-5592,-5577,-5400,-5399,-5409,-5391,-5350,-5344,-5333,-5286,-5137,-5071,-4789,-4949,-5045,-5079,-5046,-5010,-5001,-4977,-5006,-4984,-4940,-4791,-4866,-4891,-4926,-4949,
		-5498,-5506,-5499,-5511,-5521,-5558,-5474,-5023,-5496,-5595,-5338,-4703,-5473,-5488,-5572,-5604,-5607,-5606,-5600,-5588,-5566,-5549,-5549,-5550,-5572,-5601,-5603,-5594,-5598,-5599,-5680,-5589,-5636,-5461,-5400,-5398,-5394,-5304,-5299,-5298,-5230,-5130,-4658,-3057,-4930,-4975,-5004,-5010,-4997,-4968,-4972,-4978,-4952,-4799,-4781,-4789,-4830,-4912,-4953,
		-5500,-5502,-5500,-5508,-5518,-5540,-5327,-4728,-5497,-5565,-5494,-5488,-5520,-5561,-5596,-5624,-5617,-5597,-5574,-5562,-5548,-5502,-5500,-5513,-5547,-5569,-5567,-5563,-5570,-5558,-5545,-5489,-5399,-5416,-5392,-5392,-5290,-5203,-5202,-5153,-5200,-5180,-4931,-4907,-5011,-5012,-4997,-4966,-4941,-4929,-4931,-4938,-4944,-4789,-3758,-4604,-4803,-4943,-4999,
		-5445,-5497,-5504,-5506,-5513,-5523,-5539,-5519,-5557,-5578,-5553,-5565,-5572,-5585,-5602,-5607,-5588,-5555,-5542,-5539,-5527,-5506,-5498,-5498,-5512,-5530,-5540,-5542,-5539,-5518,-5499,-5444,-5393,-5401,-5358,-5211,-5199,-5164,-5159,-5159,-5191,-5181,-5173,-4955,-4947,-4990,-4901,-4865,-4850,-4897,-4895,-4888,-4816,-4871,-4778,-4784,-4829,-4946,-4995,
		-5406,-5463,-5490,-5499,-5512,-5518,-5499,-5546,-5578,-5586,-5576,-5558,-5564,-5572,-5579,-5569,-5550,-5530,-5529,-5528,-5524,-5511,-5505,-5499,-5495,-5505,-5515,-5528,-5510,-5478,-5461,-5424,-5401,-5405,-5208,-5195,-5126,-5110,-5098,-5087,-5036,-4992,-4178,-4782,-4774,-4652,-4755,-4791,-4801,-4806,-4826,-4816,-4494,-4772,-4688,-4884,-4981,-4942,-4899,
		-5402,-5432,-5474,-5495,-5500,-5500,-5518,-5548,-5570,-5586,-5577,-5563,-5561,-5562,-5561,-5552,-5537,-5501,-5501,-5529,-5526,-5514,-5508,-5499,-5492,-5496,-5499,-5515,-5492,-5453,-5433,-5405,-5397,-5421,-5206,-5125,-5065,-5083,-5075,-5060,-5002,-4991,-4575,-4766,-4572,-4447,-4765,-4791,-4803,-4801,-4802,-4814,-4565,-4589,-4233,-4826,-4887,-4834,-4806,
		-5391,-5402,-5462,-5486,-5499,-5500,-5501,-5548,-5558,-5574,-5573,-5559,-5548,-5541,-5536,-5531,-5529,-5501,-5501,-5502,-5529,-5527,-5515,-5494,-5470,-5452,-5483,-5498,-5452,-5395,-5376,-5350,-5329,-5334,-5199,-5069,-5003,-5019,-5021,-5004,-4985,-4905,-4793,-4561,-3131,-4222,-4610,-4700,-4805,-4806,-4808,-4805,-4786,-4323,-4712,-4670,-4732,-4839,-4895,
		-5407,-5422,-5467,-5497,-5500,-5500,-5501,-5522,-5537,-5553,-5555,-5539,-5526,-5523,-5520,-5520,-5529,-5501,-5516,-5530,-5527,-5523,-5501,-5476,-5428,-5401,-5403,-5402,-5351,-5307,-5283,-5234,-5188,-5187,-5186,-5072,-4999,-4940,-4998,-4998,-4951,-4935,-4739,-4477,-4701,-4746,-4749,-4760,-4780,-4804,-4801,-4799,-4791,-4605,-4786,-4785,-4797,-4805,-4987,
		-5472,-5469,-5482,-5499,-5505,-5513,-5547,-5504,-5501,-5529,-5545,-5504,-5501,-5501,-5505,-5510,-5520,-5525,-5528,-5526,-5518,-5496,-5449,-5376,-5314,-5315,-5313,-5294,-5286,-5236,-5185,-5174,-5086,-5048,-5003,-5000,-4966,-4890,-4882,-4854,-4804,-4805,-4785,-4749,-4551,-4469,-4582,-4659,-4688,-4762,-4778,-4751,-4696,-4698,-4770,-4623,-4639,-4990,-4811,
		-5500,-5497,-5497,-5499,-5503,-5515,-5523,-5546,-5501,-5502,-5523,-5500,-5495,-5495,-5498,-5500,-5507,-5511,-5516,-5498,-5471,-5395,-5345,-5302,-5275,-5261,-5255,-5249,-5231,-5191,-5164,-5059,-5000,-4950,-4942,-4946,-4946,-4824,-4758,-4712,-4600,-4684,-4587,-4458,-2610,-3960,-3968,-4290,-4593,-4703,-4739,-4670,-4609,-4617,-4809,-4904,-4995,-4808,-4956,
		-5504,-5498,-5495,-5497,-5505,-5514,-5516,-5532,-5503,-5502,-5514,-5497,-5497,-5497,-5499,-5500,-5500,-5498,-5493,-5492,-5426,-5357,-5308,-5281,-5262,-5244,-5235,-5224,-5201,-5195,-5191,-5038,-4998,-4912,-4914,-4913,-4915,-4854,-4600,-4364,-4239,-4601,-4577,-4194,-3051,-2590,-3538,-4370,-4394,-4682,-4705,-4649,-4592,-4672,-4951,-5002,-4998,-4945,-4997,
		-5477,-5496,-5490,-5493,-5513,-5515,-5485,-5478,-5541,-5542,-5507,-5501,-5501,-5503,-5502,-5497,-5478,-5441,-5406,-5383,-5364,-5322,-5302,-5274,-5250,-5231,-5206,-5202,-5159,-5172,-5168,-5014,-4953,-4877,-4852,-4856,-4907,-4751,-3065,-1281,-4371,-4492,-4411,-4480,-4339,-2331,-3516,-3836,-4008,-4579,-4631,-4572,-4734,-4872,-4995,-4954,-4901,-4888,-4976,
		-5450,-5400,-5401,-5402,-5481,-5493,-5465,-5438,-5471,-5472,-5500,-5504,-5501,-5503,-5504,-5493,-5455,-5365,-5304,-5304,-5303,-5298,-5277,-5249,-5228,-5209,-5184,-5151,-5102,-5042,-5024,-5001,-4996,-4807,-4742,-4691,-4735,-4686,-4226,-3074,-4162,-4401,-4394,-4490,-4176,-4402,-4134,-3048,-3518,-4461,-4469,-4503,-4916,-4979,-4664,-4684,-4767,-4339,-2353,
		-5490,-5458,-5404,-5398,-5401,-5406,-5334,-5117,-5065,-5492,-5512,-5511,-5503,-5500,-5501,-5498,-5478,-5354,-5278,-5271,-5264,-5250,-5238,-5213,-5196,-5170,-5147,-5118,-5077,-5006,-4991,-4996,-4977,-4803,-4239,-4396,-4581,-4489,-4550,-4350,-1859,-3657,-4134,-4391,-4500,-4577,-4303,-3631,-2600,-4408,-4373,-3707,-3075,-4767,-4306,-3061,-3502,-4211,-4192,
		-5449,-5497,-5450,-5400,-5395,-5394,-5324,-5161,-5028,-5379,-5501,-5506,-5498,-5496,-5503,-5497,-5497,-5306,-5272,-5258,-5248,-5228,-5214,-5197,-5167,-5140,-5119,-5096,-5057,-5007,-4955,-4995,-4950,-4803,-3455,-3125,-4567,-4393,-4557,-4358,-2157,-3493,-3971,-4278,-4496,-4535,-4188,-3334,-2872,-4394,-4558,-4368,-3130,-4419,-4250,-2996,-2084,-3887,-4338,
		-5161,-5152,-5494,-5451,-5209,-5087,-5392,-5395,-5395,-5403,-5442,-5456,-5485,-5497,-5522,-5536,-5547,-5370,-5216,-5222,-5225,-5197,-5179,-5150,-5116,-5082,-5056,-5049,-5024,-4980,-4854,-4798,-4868,-4818,-4416,-4170,-4364,-4005,-4467,-4465,-4354,-3252,-2709,-4100,-4484,-4518,-4219,-3067,-3976,-4430,-4576,-4478,-4114,-3966,-2652,-1424,-921,-1371,-3242,
		-5391,-5398,-5400,-5395,-5206,-5060,-5212,-5413,-5436,-5494,-5466,-5461,-5400,-5358,-5489,-5474,-5464,-5285,-5170,-5157,-5148,-5127,-5117,-5095,-5055,-5016,-4994,-4978,-4935,-4832,-4773,-4744,-4783,-4773,-4650,-4464,-4367,-2734,-4240,-4383,-4381,-4135,-3980,-3526,-4366,-4458,-4407,-4424,-3540,-4388,-4592,-4591,-4242,-3940,-1991,-0,-0,-0,-993,
		-5348,-5354,-5339,-5304,-5296,-5294,-5296,-5332,-5371,-5484,-5497,-5511,-5349,-5118,-5023,-5202,-5199,-5192,-5073,-5044,-5035,-5043,-5050,-5045,-5002,-4966,-4918,-4871,-4820,-4757,-4721,-4672,-4678,-4596,-4589,-4478,-4386,-4387,-4396,-4400,-4398,-4267,-3860,-3973,-3688,-3979,-3954,-3057,-4349,-4486,-4642,-4602,-4399,-3586,-2428,-0,-0,-0,-0,
		-5321,-5316,-5307,-5301,-5256,-5203,-5202,-5204,-5253,-5302,-5360,-5423,-5482,-5478,-5201,-5197,-5012,-4984,-4998,-5000,-4999,-5015,-5029,-5045,-5011,-4935,-4835,-4765,-4726,-4683,-4654,-4587,-4586,-4556,-4490,-4387,-4026,-4382,-4385,-4385,-4366,-4332,-3819,-3747,-3835,-3658,-3072,-3980,-2921,-4613,-4576,-4608,-4393,-3908,-1934,-0,-0,-0,-0,
		-5300,-5298,-5300,-5300,-5295,-5233,-5201,-5202,-5204,-5206,-5270,-5302,-5479,-5477,-5470,-5193,-5192,-5003,-4975,-4952,-4943,-4957,-4971,-5002,-5006,-4908,-4786,-4722,-4689,-4653,-4621,-4582,-4554,-4513,-4479,-4383,-4023,-4340,-4339,-4320,-4252,-4128,-3797,-3709,-3815,-3987,-3091,-3851,-4024,-4616,-4592,-4654,-4381,-2984,-1457,-0,-0,-0,-0,
		-5261,-5257,-5207,-5254,-5247,-5228,-5197,-5188,-5202,-5198,-5184,-5158,-5127,-5099,-5011,-5009,-5097,-5076,-4938,-4679,-4627,-4625,-4626,-4789,-4845,-4780,-4712,-4666,-4638,-4610,-4591,-4589,-4533,-4459,-4412,-4384,-4024,-4271,-4278,-4257,-4145,-3944,-3741,-3697,-3923,-4005,-4441,-4576,-4591,-4489,-4429,-4647,-4518,-2927,-0,-0,-0,-0,-0,
		-5188,-5224,-5218,-5198,-5165,-5147,-5191,-5191,-5141,-5117,-5084,-5065,-5028,-4999,-4977,-4977,-4970,-4966,-4884,-4678,-4598,-4579,-4559,-4621,-4708,-4703,-4675,-4633,-4604,-4589,-4585,-4582,-4546,-4488,-4274,-4388,-4255,-4291,-4141,-3993,-4157,-3977,-3786,-3976,-3990,-4203,-4588,-4644,-4705,-4701,-4654,-4504,-4043,-1387,-55,-0,-0,-0,-0,
		-5007,-5102,-5110,-5090,-5053,-5041,-4993,-4943,-4998,-4958,-4929,-4924,-4918,-4900,-4866,-4857,-4846,-4830,-4766,-4636,-4486,-4046,-4590,-4627,-4698,-4691,-4650,-4613,-4595,-4565,-4553,-4536,-4502,-4335,-4183,-4333,-4353,-4316,-4307,-4394,-4384,-4004,-3996,-4001,-3814,-4144,-4496,-4590,-4591,-4597,-4572,-4267,-2081,-1069,-383,-75,-0,-0,-0,
		-4990,-4986,-4996,-5002,-4971,-4981,-4982,-4882,-4913,-4887,-4848,-4803,-4801,-4794,-4786,-4782,-4766,-4755,-4725,-4645,-4501,-4320,-4594,-4668,-4691,-4673,-4639,-4605,-4584,-4556,-4542,-4517,-4485,-4353,-4267,-4363,-4385,-4321,-4395,-4399,-4394,-3839,-4134,-4378,-4016,-4024,-4392,-4566,-4310,-4271,-4123,-3946,-2070,-1062,-499,-0,-0,-0,-727,
		-4740,-4733,-4820,-4860,-4967,-4602,-4064,-4713,-4743,-4705,-4700,-4653,-4672,-4700,-4682,-4679,-4666,-4674,-4692,-4697,-4669,-4664,-4681,-4681,-4633,-4630,-4620,-4599,-4585,-4553,-4537,-4513,-4483,-4409,-4391,-4398,-4355,-4281,-4402,-4455,-4519,-4557,-4592,-4593,-4408,-4030,-4174,-4132,-2995,-2995,-3584,-2986,-2336,-1692,-509,-0,-38,-520,-1047,
		-4739,-4704,-4696,-4690,-4602,-4598,-4611,-4634,-4646,-4641,-4630,-4623,-4634,-4640,-4645,-4640,-4637,-4645,-4664,-4677,-4679,-4672,-4659,-4631,-4600,-4601,-4616,-4617,-4603,-4570,-4552,-4509,-4485,-4440,-4401,-4339,-4146,-4161,-4402,-4509,-4635,-4603,-4733,-4794,-4501,-4257,-3027,-2524,-1091,-1062,-1960,-1960,-1952,-1926,-1099,-1076,-1030,-1661,-2314,
		-4755,-4718,-4698,-4699,-4650,-4619,-4597,-4596,-4600,-4600,-4600,-4598,-4596,-4596,-4596,-4597,-4599,-4612,-4623,-4627,-4624,-4601,-4600,-4598,-4582,-4602,-4629,-4655,-4664,-4618,-4582,-4542,-4489,-4465,-4399,-4349,-4013,-4015,-4399,-4511,-4588,-4607,-4474,-4505,-4641,-4899,-2956,-1999,-919,-531,-0,-503,-515,-979,-1902,-1947,-2167,-2915,-2666,
		-4746,-4718,-4705,-4698,-4686,-4652,-4606,-4601,-4593,-4590,-4589,-4581,-4568,-4563,-4562,-4566,-4572,-4594,-4599,-4600,-4596,-4595,-4573,-4564,-4564,-4597,-4625,-4670,-4701,-4659,-4614,-4566,-4522,-4490,-4491,-4397,-4099,-4020,-4397,-4399,-4449,-4428,-3683,-3559,-3730,-4333,-2916,-1663,-532,-276,-82,-23,-0,-0,-0,-1637,-1949,-2031,-2098,
		-4724,-4716,-4709,-4706,-4702,-4702,-4684,-4633,-4591,-4585,-4577,-4549,-4507,-4491,-4485,-4495,-4512,-4531,-4544,-4543,-4527,-4499,-4474,-4464,-4472,-4525,-4598,-4649,-4764,-4735,-4679,-4581,-4547,-4565,-4582,-4589,-4315,-4181,-4379,-4007,-3670,-3016,-3567,-1737,-2628,-1993,-1921,-984,-0,-10,-0,-0,-0,-0,-452,-1466,-1858,-2702,-3981,
		-4697,-4700,-4700,-4700,-4700,-4700,-4710,-4675,-4607,-4594,-4583,-4530,-4448,-4437,-4417,-4444,-4455,-4475,-4490,-4486,-4461,-4403,-4401,-4412,-4426,-4447,-4470,-4597,-4698,-4722,-4641,-4554,-4531,-4457,-4566,-4609,-4619,-4442,-3976,-3538,-3017,-2452,-1045,-567,-547,-821,-488,-471,-72,-31,-0,-114,-362,-527,-1487,-2546,-3494,-4208,-4700,
		-4634,-4654,-4664,-4663,-4660,-4657,-4668,-4659,-4608,-4602,-4599,-4515,-4437,-4431,-4117,-4342,-4417,-4427,-4450,-4448,-4402,-4398,-4363,-4312,-4247,-4412,-4405,-4443,-4534,-4535,-4533,-4338,-4130,-3994,-4389,-4575,-4561,-4106,-3010,-2969,-2659,-556,-511,-497,-487,-311,-0,-0,-0,-0,-61,-180,-581,-1079,-2993,-4054,-4555,-4989,-5349,
		-4576,-4600,-4616,-4618,-4601,-4601,-4601,-4601,-4599,-4593,-4590,-4529,-4428,-4194,-3598,-4302,-4368,-4399,-4428,-4430,-4400,-4310,-4302,-4214,-4023,-4055,-4270,-4454,-4446,-4242,-4248,-3996,-3812,-3872,-4360,-4636,-4559,-3044,-2415,-2329,-1266,-0,-0,-0,-488,-570,-554,-721,-1050,-1071,-1093,-1124,-1620,-2588,-4015,-4978,-5121,-5387,-5472,
		-4553,-4572,-4594,-4597,-4583,-4580,-4581,-4583,-4582,-4578,-4571,-4536,-4305,-4191,-4016,-4434,-4362,-4392,-4424,-4422,-4400,-4311,-4307,-4010,-3435,-3985,-4019,-4170,-4237,-4243,-4150,-3889,-3724,-3850,-4359,-4574,-4330,-3023,-2218,-1995,-739,-0,-0,-0,-628,-731,-1069,-1995,-2486,-2667,-2552,-3042,-3529,-4459,-5062,-5157,-5357,-5399,-5400,
		-4490,-4516,-4530,-4538,-4539,-4539,-4538,-4537,-4532,-4519,-4502,-4412,-4216,-4184,-3876,-4414,-4397,-4391,-4421,-4416,-4400,-4310,-4302,-4088,-2591,-1147,-2933,-2023,-2963,-3390,-3496,-3502,-3377,-3594,-3988,-3988,-3970,-2962,-1973,-1480,-0,-0,-0,-517,-1333,-2011,-2992,-3923,-3971,-4192,-4813,-5297,-5557,-5614,-5605,-5615,-5620,-5502,-5307,
		-4415,-4444,-4469,-4487,-4490,-4489,-4484,-4480,-4474,-4458,-4434,-4394,-3944,-4186,-4129,-4396,-4411,-4393,-4408,-4400,-4393,-4349,-4291,-4156,-3006,-1601,-1975,-706,-1024,-2119,-2850,-2376,-2029,-2974,-3376,-3323,-2961,-2108,-1084,-1068,-1029,-351,-405,-1072,-2044,-3009,-3966,-4289,-4476,-4665,-5179,-5384,-5459,-5521,-5503,-5402,-5398,-5295,-5193,
		-4396,-4434,-4402,-4426,-4448,-4443,-4432,-4428,-4427,-4422,-4414,-4398,-4211,-3849,-4394,-4422,-4396,-4394,-4397,-4397,-4375,-4332,-4298,-4218,-4034,-3457,-2166,-0,-0,-839,-626,-0,-0,-722,-2406,-2948,-2064,-1932,-2082,-2988,-2984,-2517,-2375,-3313,-3809,-3973,-4227,-4302,-4296,-4975,-5087,-5197,-5297,-5309,-5204,-5196,-5192,-5001,-4809,
		-4034,-4397,-4403,-4403,-4430,-4424,-4401,-4398,-4397,-4398,-4401,-4400,-4399,-4353,-4398,-4397,-4396,-4394,-4397,-4350,-4318,-4307,-4307,-4190,-4049,-3946,-2961,-172,-391,-671,-0,-0,-0,-320,-2049,-2970,-2690,-2103,-3038,-3950,-3958,-3951,-3955,-4021,-4249,-4087,-3993,-4064,-4522,-4972,-4996,-5117,-5194,-5195,-5123,-5003,-4998,-4809,-4799,
		-4398,-4581,-4044,-4463,-4407,-4397,-4360,-4332,-4328,-4318,-4321,-4336,-4426,-4577,-4378,-4329,-4342,-4317,-4342,-4366,-4359,-4342,-4345,-4275,-4183,-4101,-3849,-2015,-2179,-849,-96,-0,-0,-0,-2039,-3405,-3956,-4103,-4493,-4567,-4658,-4767,-4766,-4771,-4595,-4580,-4110,-3571,-4278,-4108,-4788,-4820,-4810,-4809,-4805,-4798,-4713,-4679,-4603,
		-4397,-4403,-4404,-4402,-4375,-4354,-4318,-4311,-4328,-4355,-4357,-4331,-4311,-4289,-4312,-4302,-4282,-4284,-4357,-4421,-4338,-4180,-4165,-4055,-4153,-4187,-4121,-4072,-4255,-3911,-2923,-838,-1421,-1734,-2989,-3641,-4272,-4573,-4774,-4365,-4802,-4843,-4810,-4846,-4849,-4788,-4528,-4509,-4220,-4383,-4604,-4787,-4608,-4667,-4616,-4602,-4565,-4505,-4501,
		-4343,-4354,-4360,-4379,-4329,-4310,-4332,-4439,-4505,-4542,-4518,-4372,-4206,-4199,-4103,-4212,-4108,-3996,-4184,-4194,-3990,-3239,-2991,-3092,-3973,-4255,-4328,-4575,-4543,-4272,-3819,-3264,-2987,-2975,-3273,-3761,-4141,-4594,-4844,-4821,-4923,-4898,-4852,-4828,-4805,-4793,-4638,-4593,-4316,-4593,-4577,-4592,-4518,-4495,-4476,-4467,-4461,-4401,-4396,
		-4280,-4233,-4237,-4306,-4309,-4319,-4362,-4389,-4445,-4522,-4492,-4221,-3984,-3773,-3405,-3469,-3519,-3384,-3499,-3954,-3533,-1612,-281,-1440,-3041,-4183,-4323,-4738,-4668,-4507,-4267,-3903,-3858,-3766,-3832,-3993,-4213,-4785,-4786,-4819,-4865,-4818,-4796,-4796,-4713,-4684,-4599,-4593,-4474,-4497,-4492,-4406,-4389,-4391,-4323,-4342,-4335,-4296,-4265,
		-4259,-4145,-4159,-4266,-4289,-4304,-4300,-4208,-4207,-4490,-4214,-4187,-3893,-3339,-2665,-2952,-2932,-2911,-3003,-3481,-3268,-2061,-1128,-1145,-3044,-4184,-4330,-4782,-4741,-4714,-4282,-4103,-4120,-4120,-4064,-4116,-4228,-4787,-4793,-4808,-4804,-4808,-4793,-4708,-4612,-4606,-4591,-4538,-4440,-4413,-4428,-4393,-4279,-4203,-4264,-4279,-4249,-4191,-4180,
		-4180,-4240,-4164,-4188,-4175,-4175,-3971,-3798,-3933,-3929,-3845,-3376,-3046,-2927,-1085,-1059,-1953,-1977,-2035,-3184,-3465,-3933,-3918,-3301,-4006,-4234,-4486,-4827,-4817,-4840,-4922,-4230,-4372,-4555,-4517,-4516,-4592,-4662,-4772,-4787,-4732,-4686,-4654,-4599,-4577,-4504,-4461,-4447,-4396,-4390,-4385,-4199,-4144,-4107,-4099,-4167,-4162,-4051,-3988,
		-2988,-2977,-2714,-4028,-3967,-3950,-3016,-2841,-2398,-2229,-2917,-2004,-1999,-1999,-1096,-1067,-1031,-849,-1569,-3016,-3983,-4184,-4332,-4285,-4402,-4474,-4619,-4638,-4764,-4773,-4821,-4769,-4684,-4585,-4514,-4486,-4468,-4404,-4459,-4498,-4561,-4596,-4544,-4498,-4453,-4407,-4394,-4343,-4276,-4193,-4143,-4098,-4056,-4024,-4008,-3540,-3688,-3946,-3879,
		-1032,-1063,-2043,-3493,-3038,-2426,-1184,-2040,-1114,-1105,-1099,-1399,-1575,-2045,-2978,-2962,-2194,-1107,-2063,-3597,-4183,-4377,-4387,-4520,-4585,-4667,-4741,-4805,-4832,-4790,-4735,-4692,-4649,-4594,-4543,-4498,-4422,-4229,-4367,-2893,-4273,-4478,-4449,-4431,-4407,-4351,-4263,-4228,-4129,-4061,-4060,-4028,-4024,-4013,-3998,-3786,-3776,-3987,-4022,
		-534,-714,-2036,-3396,-3042,-2583,-1497,-2963,-2045,-2041,-2039,-2040,-2367,-2983,-3240,-3475,-2966,-2056,-2998,-3733,-4192,-4391,-4478,-4585,-4638,-4709,-4783,-4819,-4833,-4795,-4755,-4695,-4646,-4600,-4560,-4529,-4475,-4327,-4371,-3413,-4119,-4390,-4427,-4417,-4366,-4272,-4222,-4198,-4118,-4052,-4042,-4011,-4029,-4005,-4003,-3980,-4001,-4011,-4076,
		-429,-600,-2432,-3957,-3976,-3490,-3056,-3499,-3521,-3655,-3955,-3504,-3718,-3965,-3057,-3983,-3961,-3568,-3792,-4114,-4303,-4488,-4564,-4656,-4692,-4740,-4809,-4818,-4820,-4778,-4738,-4675,-4626,-4588,-4575,-4579,-4503,-4383,-4577,-4485,-4455,-4398,-4410,-4438,-4293,-3988,-4155,-4172,-4190,-4119,-4002,-3964,-4015,-4110,-4111,-4121,-4110,-4142,-4166,
		-542,-2010,-3484,-4284,-4375,-4195,-4189,-4005,-4096,-4256,-4382,-4388,-4387,-4387,-4391,-4310,-4194,-4189,-4193,-4294,-4402,-4546,-4609,-4690,-4710,-4792,-4812,-4802,-4787,-4735,-4696,-4631,-4580,-4524,-4544,-4574,-4560,-4518,-4519,-4589,-4590,-4400,-4411,-4394,-4231,-4104,-4075,-4104,-4179,-4174,-4088,-3970,-4104,-4192,-4196,-4189,-4186,-4190,-4199,
		-1085,-2537,-4168,-4442,-4583,-4584,-4489,-4455,-4480,-4500,-4545,-4614,-4666,-4626,-4591,-4497,-4403,-4382,-4382,-4408,-4522,-4617,-4606,-4696,-4756,-4787,-4785,-4778,-4740,-4680,-4645,-4608,-4548,-4512,-4419,-4418,-4561,-4546,-4498,-4576,-4588,-4485,-4374,-4392,-4253,-4171,-4191,-4192,-4194,-4145,-4147,-4209,-4204,-4187,-4183,-4154,-4141,-4165,-4183,
		-2104,-3963,-4436,-4622,-4641,-4636,-4653,-4655,-4691,-4709,-4756,-4926,-4661,-4593,-4419,-4581,-4538,-4446,-4504,-4567,-4604,-4695,-4656,-4632,-4709,-4769,-4763,-4752,-4690,-4624,-4601,-4567,-4563,-4570,-4581,-4566,-4560,-4472,-4586,-4582,-4389,-4348,-4271,-4211,-4329,-4388,-4225,-4081,-4143,-4197,-4206,-4102,-4086,-3934,-4201,-4164,-4125,-4155,-4202,
		-3057,-4056,-4582,-4693,-4702,-4706,-4658,-4641,-4684,-4713,-4768,-4962,-4724,-4057,-4431,-4595,-4589,-4162,-4585,-4593,-4652,-4626,-4608,-4556,-4663,-4756,-4756,-4737,-4677,-4600,-4588,-4589,-4563,-4552,-4567,-4577,-4535,-4533,-4587,-4425,-4221,-4223,-4299,-4391,-4351,-4391,-4387,-4386,-4235,-4293,-4390,-4330,-4388,-4176,-4114,-4200,-4200,-4202,-4239,
		-4575,-4561,-4699,-4830,-4891,-4904,-4884,-4994,-4851,-4759,-4705,-4699,-4710,-4630,-4617,-4569,-4456,-4460,-4346,-4614,-4674,-4452,-4407,-4045,-4313,-4732,-4768,-4697,-4619,-4544,-4541,-4577,-4622,-4616,-4571,-4603,-4580,-4560,-4592,-4501,-4406,-4398,-4215,-4393,-4394,-4396,-4288,-4396,-4398,-4398,-4398,-4288,-4395,-4393,-4402,-4329,-4297,-4397,-4400,
		-4845,-4746,-4893,-4964,-4992,-4996,-5000,-5014,-4974,-4848,-4759,-4723,-4701,-4702,-4697,-4680,-4594,-4595,-4599,-4604,-4638,-4573,-4566,-4279,-4616,-4823,-4842,-4835,-4754,-4254,-4412,-4512,-4546,-4551,-4534,-4545,-4557,-4560,-4570,-4590,-4586,-4570,-4538,-4497,-4336,-4438,-4483,-4480,-4472,-4446,-4404,-4390,-4390,-4334,-4381,-4372,-4386,-4433,-4383,
		-4982,-4970,-4999,-5020,-5028,-5017,-5004,-4996,-4930,-4840,-4797,-4788,-4787,-4790,-4804,-4797,-4773,-4704,-4700,-4690,-4592,-4573,-4385,-4173,-4606,-4735,-4793,-4718,-4595,-4538,-4529,-4559,-4573,-4570,-4551,-4573,-4452,-4556,-4575,-4584,-4596,-4590,-4593,-4587,-4544,-4594,-4587,-4588,-4562,-4577,-4216,-4398,-4377,-4402,-4403,-4439,-4465,-4589,-4506,
		-4997,-4998,-5012,-5021,-5025,-5019,-4998,-4987,-4892,-4829,-4802,-4810,-4821,-4824,-4834,-4865,-4798,-4755,-4720,-4645,-4569,-4576,-4570,-4342,-4524,-4672,-4726,-4701,-4619,-4586,-4585,-4592,-4598,-4590,-4547,-4433,-4420,-4562,-4577,-4578,-4583,-4544,-4591,-4382,-4586,-4595,-4595,-4590,-4575,-4571,-4104,-4509,-4476,-4408,-4425,-4394,-4462,-4602,-4604,
		-4982,-4974,-4970,-4968,-4964,-4957,-4915,-4866,-4833,-4815,-4807,-4808,-4818,-4811,-4782,-4672,-4740,-4780,-4773,-4649,-4596,-4588,-4585,-4581,-4347,-4542,-4678,-4725,-4611,-4544,-4560,-4639,-4606,-4606,-4520,-4483,-4473,-4582,-4640,-4618,-4601,-4601,-4560,-4582,-4586,-4545,-4420,-4096,-3784,-4577,-4498,-4477,-4614,-4631,-4594,-4590,-4592,-4609,-4703,
			;
}
